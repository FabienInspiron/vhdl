library IEEE;
use IEEE.numeric_bit.all;

architecture archi_decoder of decoder is
	
begin
		
				
end architecture archi_decoder;
