ENTITY testbench IS
END testbench;